`include "riscv/src/defines.v"

module RegFile(
    input wire clk,
    input wire rst,
    input wire rdy

);


endmodule