`include "riscv/src/defines.v"

module InstFetcher(
    input wire clk,
    input wire rst,
    input wire rdy

    
);

endmodule