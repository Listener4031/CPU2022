module ALUnit();

endmodule