`include "riscv/src/defines.v"

module InstCache(
    input wire clk,
    input wire rst,
    input wire rdy

    // InstFetcher

    // MemController
);

endmodule