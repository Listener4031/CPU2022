module Test(
    input wire clk,
    input wire rst
);



endmodule