module LSBuffer(
    input wire clk,
    input wire rst,
    input wire rdy

    // Decoder

    // ALU_LS

    // ReorderBuffer

);

endmodule