module RegFile(
    input wire clk,
    input wire rst,
    input wire rdy,
    input wire clear
);



endmodule