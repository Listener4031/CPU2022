module CPU(
    input wire clock_in,
    input wire reset_in,
    input wire ready_in

    
);



endmodule