module ReorderBuffer(
    input wire clk,
    input wire rst,
    input wire rdy

    // Decoder
    
);

endmodule