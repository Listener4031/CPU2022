module Dispatcher(
    input wire clk,
    input wire rst,
    input wire rdy

    //Fetcher

    //ReorderBuffer

    //RegFile

    //RsvStation

    //LSBuffer

    //CDB
);

endmodule