module LSUnit();

endmodule